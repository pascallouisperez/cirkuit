innerBorder = 248,137,275,157,299,170,320,177,339,180,359,179,380,175,400,170,419,167,435,168,446,177,452,194,455,218,459,246,466,275,479,302,501,324,529,343,560,357,590,368,616,377,635,384,642,389,648,394,639,397,619,400,587,403,548,406,507,410,469,415,438,421,419,429,403,439,392,448,381,460,367,475,352,494,341,516,353,530,377,532,456,523,561,507,672,486,774,463,849,439,884,417,886,399,864,383,830,371,794,362,764,357,741,354,724,352,709,348,696,340,683,327,671,311,661,291,654,270,650,249,651,229,655,210,661,192,669,174,676,157,683,141,693,129,710,126,738,136,781,163,841,210,911,270,982,337,1045,402,1091,459,1113,501,1119,529,1122,551,1120,565,1114,598,1102,613,1058,623,894,660,684,703,462,744,261,776,116,792,77,783,68,758,94,737,148,712,192,685,189,663,173,639,140,603,115,571,92,491,79,391,74,287,79,192,94,121,118,84,148,76,182,89,216,112
tolerance = 10
name = Bahrain
maximumSpeed = 12
startingLine = 539,791,539,724
outerBorder = 97,700,53,730,15,755,6,782,13,809,43,832,205,829,426,800,671,760,904,715,1088,673,1142,658,1167,630,1177,597,1180,571,1182,552,1184,535,1186,511,1179,477,1154,430,1104,368,1034,297,955,225,876,160,806,109,752,78,714,66,686,69,666,83,650,105,635,132,620,161,609,193,602,226,600,258,609,286,619,311,635,334,654,356,668,368,685,386,704,394,724,397,742,398,762,400,783,403,795,408,789,416,760,427,702,442,626,459,543,476,467,490,410,500,395,501,387,495,397,484,415,470,433,466,468,460,515,452,565,442,613,431,651,420,673,408,681,396,677,384,664,371,646,359,625,347,602,333,580,317,560,297,543,271,530,239,520,203,511,168,500,137,485,115,465,104,441,102,416,105,391,111,368,117,349,119,332,116,312,108,287,93,254,70,210,41,160,14,110,0,64,10,28,54,7,139,0,251,6,374,24,490,51,582,85,638,107,656,134,678
