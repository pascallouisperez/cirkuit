innerBorder = 499,129,537,157,527,229,513,250,464,238,403,222,373,268,404,297,465,324,382,371,415,492,380,521,358,431,304,483,324,420,313,323,262,318,246,402,224,441,188,441,149,425,113,366,117,336,139,302,177,277,198,271,215,259,229,232,226,206,206,190,154,174,122,167,106,136,110,113,143,91,207,127,269,158,332,131,283,63,363,65,397,122,440,151
tolerance = 10
name = Complex
maximumSpeed = 7
startingLine = 144,392,144,520
outerBorder = 491,77,562,96,580,149,583,238,538,290,440,264,496,304,453,396,460,449,449,512,397,550,326,557,343,485,271,545,280,393,268,463,243,495,193,498,139,485,93,452,64,408,53,362,64,325,91,295,121,270,165,252,177,236,168,218,144,213,79,199,61,182,44,158,33,123,38,94,61,56,116,34,177,46,281,123,237,63,257,25,358,10,416,36,452,102
