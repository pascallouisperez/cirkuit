innerBorder = 201,52,249,54,303,57,357,60,407,64,448,69,476,75,494,81,503,88,506,95,507,102,507,109,507,116,506,123,502,130,496,138,487,146,475,154,462,160,449,165,436,166,424,164,414,159,404,153,394,147,384,143,374,141,364,142,355,145,347,150,341,156,338,163,336,172,336,181,337,191,338,201,338,212,339,222,340,232,343,241,348,249,356,255,365,259,376,261,387,262,398,260,408,256,416,251,425,246,434,241,444,238,455,237,467,239,480,243,492,250,503,260,513,273,520,289,524,306,524,324,517,343,504,361,486,376,466,385,445,386,425,376,408,354,395,326,383,301,372,287,361,292,350,322,341,368,336,422,339,472,351,508,374,523,404,522,434,512,458,502,472,500,470,511,455,533,431,559,402,584,371,602,343,609,318,604,299,587,285,558,279,516,280,463,287,407,294,354,300,315,299,296,290,304,273,330,249,366,221,399,190,420,158,421,129,406,108,381,100,353,110,328,140,311,181,300,223,294,254,289,263,283,243,274,204,262,160,250,122,237,106,226,120,217,155,211,197,205,233,199,250,191,238,181,205,170,163,158,125,146,101,136,81,97,83,68,117,49,134,49,162,50
tolerance = 10
name = Treesy
maximumSpeed = 10
startingLine = 461,81,461,11
outerBorder = 13,53,20,39,44,26,81,15,128,6,183,1,243,0,303,2,362,7,415,14,459,21,491,28,513,36,527,45,536,56,541,69,545,84,549,101,552,118,555,134,559,147,563,157,565,163,563,169,553,174,534,180,504,188,395,206,531,190,555,214,571,249,578,289,578,329,571,363,559,388,542,404,523,414,504,420,486,424,470,428,457,431,445,431,434,429,424,423,413,412,389,371,403,405,405,419,403,431,400,441,397,448,398,453,405,455,420,454,441,452,465,449,488,449,508,452,521,460,528,472,529,490,524,512,513,538,497,568,475,599,448,627,416,648,378,659,335,657,292,644,252,620,221,589,202,551,256,417,194,547,156,525,114,481,72,426,36,371,11,326,0,299,1,288,14,288,35,292,62,297,93,297,124,294,151,290,170,285,177,283,169,284,149,286,122,289,93,289,67,284,47,274,34,259,26,242,23,225,23,211,26,201,32,195,41,191,54,189,72,188,94,187,155,189,92,188,66,178,43,161,24,140,12,119,8,99
