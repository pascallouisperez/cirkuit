innerBorder = 491,147,496,154,501,162,506,171,511,181,515,189,518,196,519,203,521,209,522,214,523,219,525,224,527,229,528,234,528,239,527,243,524,246,519,249,513,250,506,251,498,250,490,248,482,246,473,242,464,238,454,234,443,230,432,226,422,223,412,221,403,222,396,225,390,231,385,239,381,248,377,258,373,268,370,279,369,287,371,294,378,298,389,298,404,297,420,294,436,294,450,296,460,303,465,313,465,324,461,334,451,343,436,348,418,350,399,349,381,347,366,344,356,341,352,341,350,344,352,354,355,372,359,399,363,432,366,465,368,494,368,514,366,521,361,518,356,509,351,496,346,483,343,473,340,467,339,462,338,459,337,456,336,453,335,449,333,445,332,440,330,434,328,428,327,421,325,415,324,409,322,403,320,398,318,394,316,390,312,386,306,381,299,375,290,370,281,364,272,361,265,359,259,360,255,364,253,370,251,377,249,385,247,393,246,402,244,410,241,418,238,425,234,431,229,437,224,441,218,443,212,445,206,445,200,444,194,443,188,441,182,439,176,438,170,436,163,434,156,431,149,425,141,417,134,407,127,396,121,385,116,375,113,366,112,359,112,354,113,348,114,344,115,340,117,336,118,331,121,326,124,321,128,315,133,308,139,302,145,295,152,290,159,286,165,282,171,279,177,277,182,276,186,275,190,274,193,273,195,272,198,271,201,269,203,268,206,265,209,263,212,261,215,259,218,256,221,253,224,250,226,245,228,239,229,232,230,225,230,219,230,214,229,210,228,208,226,206,224,205,222,203,219,200,216,197,211,193,206,190,199,186,191,183,181,180,172,177,162,175,154,174,147,173,141,173,136,173,131,172,127,170,122,167,118,163,114,158,110,153,108,147,107,142,106,136,107,131,107,127,108,123,108,120,109,116,110,113,112,110,115,107,120,103,127,99,135,95,143,91,152,88,160,85,168,83,175,81,182,80,187,78,191,76,195,75,199,74,203,72,209,71,217,70,226,69,236,69,247,68,257,68,267,68,275,68,283,68,290,68,297,68,303,68,309,69,314,69,321,71,328,72,337,74,346,76,356,79,366,81,375,84,384,87,392,89,400,92,408,96,417,100,427,105,437,111,448,117,458,122,466,127,473,131,478,134,482,138,487,142
tolerance = 10
name = Complex
maximumSpeed = 9
startingLine = 144,100,30,100
outerBorder = 487,43,501,51,516,60,530,70,543,80,554,89,562,96,567,103,571,109,574,116,576,125,578,136,580,149,582,163,584,179,585,194,585,209,585,224,583,238,580,250,576,262,570,272,562,280,551,286,538,290,521,290,501,287,481,283,462,276,448,270,440,264,441,260,449,259,461,261,474,269,487,283,496,304,501,328,502,353,497,375,487,390,472,396,453,396,434,393,416,389,403,390,396,397,395,409,397,425,401,442,405,459,408,474,409,487,410,499,409,509,407,519,404,528,401,536,396,543,390,548,382,551,373,551,362,549,352,546,343,542,335,538,330,534,326,531,324,528,322,524,320,520,317,515,314,509,310,504,307,499,304,495,302,492,300,490,298,486,296,481,294,471,291,457,288,441,285,425,282,414,279,408,277,411,274,420,272,434,270,449,268,463,265,474,262,481,258,487,254,490,249,493,243,495,237,497,230,499,222,500,213,500,203,499,193,498,183,496,173,494,163,492,154,490,146,487,139,485,132,481,124,477,116,472,108,466,100,459,93,452,86,445,80,438,75,430,71,423,67,416,64,408,61,400,58,392,56,384,54,377,53,369,53,362,54,355,55,348,57,342,59,336,61,330,64,325,66,319,70,314,74,309,79,304,85,299,91,295,97,290,103,286,108,282,113,277,117,274,121,270,124,267,127,264,130,262,132,261,134,259,136,257,138,255,139,253,141,250,144,247,148,244,153,241,159,237,164,234,168,230,169,228,167,226,162,225,155,224,147,224,139,223,132,222,125,221,118,219,112,217,105,214,98,211,91,207,85,203,79,199,74,195,70,192,67,189,65,187,63,185,61,182,59,179,56,176,53,172,50,168,47,163,44,158,41,152,39,146,37,140,35,134,34,128,33,123,33,118,33,113,34,108,35,103,36,99,38,94,40,89,43,83,46,76,50,69,55,62,61,56,68,50,77,45,86,42,96,39,106,36,116,34,125,32,133,29,140,27,149,24,158,22,169,20,180,17,192,15,205,13,218,12,231,11,243,11,255,11,267,11,279,11,291,11,303,11,314,11,325,11,336,11,346,11,355,12,364,13,373,14,382,15,391,17,400,19,409,21,418,23,428,25,438,27,449,29,461,33,473,37
