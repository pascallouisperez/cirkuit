innerBorder = 328,116,349,141,351,168,335,215,367,232,367,283,347,326,333,348,365,379,380,416,375,467,368,483,347,485,336,474,322,431,310,400,290,367,264,344,174,334,258,335,311,329,337,315,353,297,356,276,354,257,347,243,332,231,319,221,177,221,288,218,323,206,329,191,335,169,334,149,320,129,292,120,115,107,291,107
tolerance = 10
name = Mega Curvy
maximumSpeed = 7
startingLine = 359,260,453,260
outerBorder = 416,144,424,192,441,235,441,284,397,341,434,361,456,401,458,443,430,498,388,529,342,539,289,529,262,505,242,459,225,426,190,408,147,406,106,414,72,395,53,366,48,327,55,306,68,292,132,282,282,272,130,276,93,273,65,267,47,251,39,226,53,200,70,183,100,168,286,163,98,160,55,149,35,117,42,89,82,64,127,55,196,51,272,53,360,71,405,113
