innerBorder = 186,231,189,248,194,263,201,274,209,282,220,289,233,294,247,297,264,299,283,299,305,299,329,298,353,295,374,288,390,278,398,262,396,240,387,214,377,187,369,161,367,139,375,123,391,114,409,113,428,118,442,132,449,153,449,180,443,209,434,239,421,267,407,290,395,310,387,325,388,336,400,344,425,349,459,352,496,355,531,358,559,362,575,369,583,377,587,388,592,400,602,412,619,425,637,437,646,450,637,463,600,475,531,487,440,497,345,506,260,512,201,514,180,513,190,508,220,500,259,489,295,477,320,463,334,449,340,434,341,420,340,406,339,393,337,381,333,370,327,360,317,351,303,343,284,335,263,328,240,323,216,319,192,316,169,315,150,314,136,313,129,311,130,308,136,304,147,295,159,283,170,265,178,241,183,215,186,189,187,170,187,159,186,160,185,172,184,190,185,210
tolerance = 10
name = New
maximumSpeed = 9
startingLine = 413,575,413,494
outerBorder = 130,147,131,130,134,112,141,96,150,81,163,71,179,65,198,63,217,65,234,69,248,76,257,84,262,93,262,104,260,116,256,129,250,143,244,158,238,173,233,186,229,199,228,210,229,219,232,226,239,232,249,236,262,239,277,242,293,244,308,245,321,246,331,247,338,245,341,241,341,231,336,215,328,191,318,163,310,133,305,106,308,85,319,72,339,67,364,67,395,70,429,73,465,76,499,78,528,81,551,85,562,93,561,104,550,120,533,138,514,159,497,183,486,208,480,234,482,257,489,275,504,286,525,289,550,287,578,284,604,284,627,290,645,306,658,329,667,357,675,386,681,412,687,434,692,451,693,466,689,480,679,493,661,507,636,522,607,535,576,547,546,556,517,561,489,563,459,564,425,564,385,565,338,567,286,570,234,572,186,571,145,566,115,556,96,543,87,527,86,511,94,496,109,484,128,473,150,464,173,456,194,447,212,437,225,427,234,415,239,404,240,391,236,378,229,366,218,357,206,351,193,349,180,353,166,360,151,369,135,375,118,378,99,375,80,366,63,354,49,339,41,322,40,305,45,289,54,274,66,260,80,249,94,240,106,233,117,226,126,220,132,212,134,203,134,191,133,178,131,163
