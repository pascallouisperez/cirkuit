innerBorder = 515,238,528,206,563,168,620,127,543,178,489,193,440,190,398,174,366,152,344,133,334,123,337,129,347,148,358,177,365,214,360,253,340,292,311,328,281,357,258,377,250,385,264,379,295,363,336,345,382,328,426,321,462,326,490,341,513,374,496,337,498,314,515,293,550,278,595,268,672,257,572,267,533,258
tolerance = 10
name = Starry
maximumSpeed = 8
startingLine = 454,100,454,204
outerBorder = 311,247,274,308,217,366,157,417,108,455,88,473,107,468,158,448,231,422,315,399,398,390,472,400,532,424,577,453,605,476,613,486,602,475,580,448,560,410,554,369,573,330,624,299,695,276,769,260,828,250,856,244,841,241,794,239,734,232,679,219,646,195,647,159,674,116,711,75,743,43,757,27,741,33,698,54,636,81,563,107,486,121,412,118,346,103,292,83,256,66,242,61,252,72,276,100,302,140,318,190
