innerBorder = 113,151,111,164,110,175,111,186,112,194,115,200,120,204,126,206,135,207,146,208,159,209,175,211,192,216,209,222,223,232,233,246,238,264,233,325,228,342,224,354,220,363,214,368,207,372,196,375,182,378,165,382,147,385,131,389,117,392,108,395,103,397,102,400,106,404,115,409,128,415,144,422,162,430,180,437,199,443,216,448,233,451,250,453,267,454,286,454,307,454,328,453,350,453,370,452,388,451,403,450,415,449,425,448,433,447,441,445,448,443,455,442,461,442,467,443,472,447,476,454,480,463,484,474,489,485,495,495,503,504,512,511,522,515,531,515,540,511,547,502,553,489,557,474,559,458,560,443,559,430,556,418,551,408,544,400,535,393,524,387,511,382,499,379,486,378,475,379,466,383,459,388,453,395,449,402,446,409,443,415,440,420,434,424,424,428,408,432,386,436,360,440,333,442,307,444,286,444,272,442,264,438,259,432,258,423,256,413,254,401,250,387,246,371,242,354,239,336,236,317,238,285,244,251,253,240,265,232,280,226,299,221,321,216,346,211,373,206,399,201,421,195,438,188,447,180,449,172,444,163,434,153,419,144,400,135,378,126,355,118,332,110,311,103,293,96,277,90,262,85,248,81,232,78,214,77,196,77,177,79,160,83,145,90,134,99,125,111,120,124,116,138
tolerance = 10
name = Big Girl
maximumSpeed = 8
startingLine = 124,187,41,187
outerBorder = 47,161,45,183,43,202,42,219,43,233,48,243,57,249,69,251,85,252,101,251,118,250,134,250,150,251,164,254,176,260,186,267,193,277,197,288,197,300,193,312,184,322,170,330,152,335,133,338,114,340,98,341,86,341,78,341,73,341,69,343,66,346,63,351,60,358,56,367,53,377,51,389,49,402,48,414,49,427,51,438,55,448,61,456,69,461,80,466,92,470,106,474,122,479,139,484,157,488,174,493,191,496,207,498,221,499,236,500,250,500,266,499,283,498,301,497,319,496,337,494,355,492,372,489,387,486,400,483,411,480,419,478,425,477,428,478,430,481,432,486,435,494,439,504,444,516,449,529,456,543,463,555,470,566,478,575,486,582,495,587,505,590,516,590,527,588,538,585,550,580,560,574,569,568,578,560,585,552,592,542,597,530,601,516,605,501,607,484,609,467,609,450,608,433,606,416,602,400,597,385,589,371,579,358,567,346,553,336,536,329,518,323,498,320,477,320,456,323,435,330,415,341,397,356,380,372,365,387,350,397,335,399,320,392,307,377,296,357,289,336,288,316,293,300,303,288,317,279,334,272,352,266,370,261,387,257,405,254,422,251,439,249,456,248,472,245,488,241,502,233,514,219,523,199,528,175,527,150,518,125,498,103,467,86,429,74,389,65,350,59,318,53,296,47,281,42,270,37,257,34,238,31,211,30,178,32,144,36,111,44,84,56,66,72,55,92,50,115,48,138
