innerBorder = 217,95,275,110,319,120,331,153,335,191,331,236,292,295,265,316,230,320,193,316,173,288,167,272,186,236,219,208,232,185,269,116
tolerance = 10
name = Patatoid
maximumSpeed = 6
startingLine = 226,236,100,236
outerBorder = 323,44,363,76,399,79,427,93,445,126,447,185,442,245,369,324,301,356,227,357,175,355,141,320,117,289,122,254,154,148,217,158,154,141,182,71,225,41,279,32
