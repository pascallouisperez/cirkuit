innerBorder = 152,180,162,172,174,162,185,152,195,142,203,132,208,122,210,113,211,105,212,97,213,90,215,84,220,78,225,74,233,71,243,70,255,71,269,73,283,76,299,80,315,84,331,88,346,93,360,97,374,102,386,106,397,111,407,116,417,121,428,128,441,135,456,144,472,152,489,160,507,166,523,168,538,166,552,160,565,150,578,136,585,114,591,92,602,71,632,58,668,49,703,39,746,35,794,37,843,43,886,51,919,60,939,69,947,78,947,86,942,94,936,102,931,110,927,117,923,124,920,131,915,138,909,144,902,150,894,156,887,161,879,165,872,169,866,172,861,174,856,177,853,180,851,183,849,187,848,192,848,199,847,207,846,217,845,229,843,242,842,255,840,268,839,280,838,290,838,300,839,309,841,318,845,326,850,334,856,340,863,345,870,348,877,349,883,348,889,345,895,342,900,337,905,332,910,327,916,323,921,320,928,321,935,325,943,331,949,340,953,349,954,359,951,369,946,378,938,387,928,396,918,405,908,414,898,424,888,433,878,442,867,450,856,457,844,464,831,470,817,475,802,480,786,484,769,488,751,491,733,494,715,498,697,502,680,506,662,508,645,508,627,505,609,498,591,490,574,481,559,474,545,472,534,475,525,483,517,492,510,502,504,510,498,514,492,515,487,513,483,509,480,503,479,497,479,490,477,482,473,475,465,469,452,463,436,458,418,453,401,447,387,440,377,432,369,424,363,415,355,407,345,401,330,397,313,394,293,393,272,393,252,395,234,398,218,401,205,405,195,409,188,414,184,419,184,424,186,429,190,435,195,441,201,447,208,454,214,463,218,473,220,486,219,501,214,518,208,535,199,549,189,561,178,568,166,572,155,573,145,573,136,573,130,574,126,576,124,579,124,584,126,591,129,600,133,609,137,619,141,628,143,635,143,640,141,642,138,642,133,642,128,641,122,640,116,639,109,638,102,636,95,634,88,631,82,628,75,624,70,618,64,611,59,602,54,592,50,580,47,566,45,551,44,535,43,518,43,500,44,482,45,464,47,447,48,430,50,415,51,400,51,386,51,373,50,361,50,348,53,334,58,318,67,299,78,279,90,259,103,240,114,224,123,211,130,202,137,194,144,187
tolerance = 10
name = Monte Carlo
maximumSpeed = 10
startingLine = 59,403,0,403
outerBorder = 7,606,13,627,20,644,30,658,41,668,54,675,69,679,84,679,100,678,116,675,131,672,145,669,156,665,166,661,173,657,178,653,180,648,179,643,177,637,174,631,172,624,171,617,170,609,171,603,173,598,176,596,180,597,186,599,191,602,198,604,204,603,210,599,216,592,221,583,225,573,229,563,232,554,234,546,237,538,239,530,243,522,248,513,253,504,257,494,260,484,260,474,257,464,252,455,247,447,241,441,238,436,237,433,240,432,244,431,252,431,261,431,272,430,285,429,298,429,311,429,323,432,334,437,343,444,353,452,363,460,375,467,389,473,403,478,417,482,429,486,438,492,443,499,445,507,446,515,449,524,454,532,463,539,476,545,490,550,503,551,515,550,524,546,530,539,534,532,538,526,543,523,549,523,557,527,567,532,579,539,593,545,609,550,626,554,645,557,665,558,685,558,706,557,727,554,748,551,769,547,789,543,809,538,827,533,845,528,861,522,876,516,889,509,901,502,911,495,921,487,929,478,937,469,944,460,950,450,957,440,963,429,969,418,975,407,981,396,986,384,991,372,995,360,998,348,999,337,999,325,996,315,991,306,984,297,975,290,966,284,957,279,948,276,939,274,931,273,923,274,915,277,907,281,900,286,893,292,887,297,882,301,878,304,876,305,875,304,874,302,875,297,876,290,878,282,880,272,882,262,884,251,885,240,887,230,889,220,892,211,897,203,904,196,914,190,924,185,935,179,945,174,954,168,962,162,969,155,975,149,979,143,982,137,984,132,986,126,986,120,986,114,986,107,985,99,983,89,980,78,976,66,970,52,961,38,944,24,919,12,883,3,808,0,718,0,663,5,618,12,587,21,568,31,558,43,554,57,553,72,551,88,548,104,542,118,532,126,517,128,497,122,473,109,448,93,424,77,402,62,385,51,371,45,359,41,347,38,332,36,314,34,294,32,272,30,251,29,231,30,214,33,199,38,187,44,178,53,172,63,168,75,166,88,164,101,161,114,156,126,147,137,136,147,122,157,107,169,91,184,75,202,59,221,45,241,32,260,21,276,13,288,7,298,3,307,1,318,0,333,0,368,0,405,0,435,0,466,0,497,0,527,1,556,3,582
