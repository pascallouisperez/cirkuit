innerBorder = 165,326,172,340,180,356,187,372,193,388,197,401,199,415,199,429,196,447,191,468,184,489,175,506,165,519,153,527,140,535,127,545,114,559,103,574,97,586,97,590,104,585,116,574,128,561,139,550,145,544,150,539,156,535,162,530,170,524,180,519,190,514,200,511,210,510,220,509,228,508,236,506,244,506,253,507,266,510,281,517,297,524,312,532,326,539,338,544,348,547,356,549,363,549,369,548,374,546,379,543,384,541,388,539,391,537,393,535,393,532,391,528,388,523,383,518,376,510,369,502,361,492,354,481,347,468,343,456,341,443,341,430,344,418,348,407,353,397,358,388,364,380,370,373,377,366,383,361,391,357,400,354,411,352,423,352,431,352,434,352,431,352,422,350,409,345,394,336,379,324,365,310,354,296,348,285,346,276,346,267,346,257,345,245,345,230,345,216,348,203,354,191,361,181,368,172,375,164,381,155,386,148,392,141,398,136,405,132,411,128,417,124,421,118,424,111,426,104,426,96,425,88,423,80,419,73,413,65,406,59,397,53,387,49,376,46,364,45,353,45,342,47,333,50,324,54,317,59,310,66,305,74,301,84,298,94,298,104,300,114,302,124,302,135,297,147,289,159,278,170,266,181,254,190,242,197,230,202,219,205,210,206,200,205,191,203,182,199,173,194,164,188,155,183,147,179,139,175,132,169,127,161,123,149,120,135,117,120,113,107,108,97,103,90,97,86,91,84,86,84,82,86,78,89,75,93,73,99,71,106,69,115,67,126,64,139,63,152,62,164,62,174,64,183,66,191,68,199,71,208,75,217,80,227,85,236,92,246,100,255,109,264,118,272,127,280,136,288,144,295,150,302,156,310,162,320
tolerance = 10
name = Biggy Curve
maximumSpeed = 8
startingLine = 2,179,70,179
outerBorder = 9,382,30,426,58,452,86,467,107,476,117,483,119,490,116,495,112,501,107,506,101,514,92,523,82,536,69,551,57,566,47,579,41,588,39,595,39,600,40,605,43,612,46,619,50,625,56,629,63,631,73,629,87,625,105,616,125,606,146,595,166,588,183,585,197,586,211,588,225,589,240,590,257,590,274,592,292,597,309,604,327,612,344,616,363,617,381,613,398,606,414,599,427,593,438,586,447,580,454,573,459,565,462,556,463,546,462,536,460,526,455,517,450,510,445,503,439,498,433,492,427,485,421,475,416,464,412,452,411,441,411,432,414,424,418,417,423,411,428,404,435,398,442,393,450,389,459,385,468,381,477,376,486,371,493,364,498,357,500,349,499,340,495,332,488,325,480,321,470,319,460,318,449,316,440,312,431,306,422,299,414,292,406,286,399,279,393,272,389,264,389,254,390,244,393,234,397,225,402,218,408,212,416,209,425,206,436,204,446,201,455,195,461,185,464,173,467,159,468,147,471,137,473,128,474,117,476,104,476,89,474,73,470,57,464,43,454,31,444,22,434,15,425,10,415,7,405,5,393,4,378,2,361,0,343,0,325,2,309,7,293,13,280,22,269,32,260,43,253,56,248,69,244,82,241,95,239,107,236,117,234,125,231,132,227,137,223,143,217,147,210,151,203,153,195,153,187,151,180,147,174,143,170,138,167,131,164,122,161,111,158,96,154,81,151,66,148,55,145,47,142,41,139,35,134,29,128,23,122,17,114,13,106,11,97,12,89,13,80,16,71,18,61,21,52,24,44,28,36,34,28,41,21,50,16,62,10,135,5,191,0,263,1,335
